-- Maquina de Vendas (Bloco Operacional)

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity BO is
	generic(
		nbits   :   integer := 8								  -- número de bits
	);
	-- Definndo as portas de entrada e saida
	port(
		clk
	);
end BO

architecture comportamento of BO is
	-- Região de declaração
	
begin -- Descrição do sistema

end architecture;